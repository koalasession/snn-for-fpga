
LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
USE ieee.std_logic_unsigned.ALL;
USE ieee.numeric_std.ALL;

ENTITY RAM_0 IS

    GENERIC (
        number : IN INTEGER;
        weight_width : IN INTEGER;
        neuron_adr : IN INTEGER;
        weights : IN INTEGER);

    PORT (
        CLK : IN STD_LOGIC;
        we : IN STD_LOGIC;
        a : IN STD_LOGIC_VECTOR(neuron_adr DOWNTO 0);
        dpra : IN STD_LOGIC_VECTOR(neuron_adr DOWNTO 0);
        di : IN STD_LOGIC_VECTOR(weights DOWNTO 0);
        dpo : OUT STD_LOGIC_VECTOR(weights DOWNTO 0));
END RAM_0;
ARCHITECTURE syn OF RAM_0 IS

    TYPE ram_type IS ARRAY (0 TO 127) OF STD_LOGIC_VECTOR(weights DOWNTO 0);
    SIGNAL RAM : ram_type := (OTHERS => (OTHERS => '0')); -- Initializes all weights to 0

BEGIN
    PROCESS (clk)
    BEGIN
        IF (rising_edge(clk)) THEN

            -- Hardcoding the weights for each neuron

            IF (number = 2) THEN

                RAM(8) <= STD_LOGIC_VECTOR(to_signed(20, RAM(19)'LENGTH));
                RAM(21) <= STD_LOGIC_VECTOR(to_signed(20, RAM(19)'LENGTH));
                RAM(39) <= STD_LOGIC_VECTOR(to_signed(20, RAM(19)'LENGTH));
                RAM(53) <= STD_LOGIC_VECTOR(to_signed(20, RAM(19)'LENGTH));
                RAM(67) <= STD_LOGIC_VECTOR(to_signed(-60, RAM(19)'LENGTH));
            ELSIF (number = 3) THEN
                RAM(43) <= STD_LOGIC_VECTOR(to_signed(20, RAM(19)'LENGTH));
                RAM(45) <= STD_LOGIC_VECTOR(to_signed(20, RAM(19)'LENGTH));
                RAM(46) <= STD_LOGIC_VECTOR(to_signed(20, RAM(19)'LENGTH));
                RAM(49) <= STD_LOGIC_VECTOR(to_signed(20, RAM(19)'LENGTH));
                RAM(65) <= STD_LOGIC_VECTOR(to_signed(-60, RAM(19)'LENGTH));
            ELSIF (number = 4) THEN
                RAM(5) <= STD_LOGIC_VECTOR(to_signed(20, RAM(19)'LENGTH));
                RAM(8) <= STD_LOGIC_VECTOR(to_signed(20, RAM(19)'LENGTH));
                RAM(12) <= STD_LOGIC_VECTOR(to_signed(20, RAM(19)'LENGTH));
                RAM(16) <= STD_LOGIC_VECTOR(to_signed(20, RAM(19)'LENGTH));
                RAM(76) <= STD_LOGIC_VECTOR(to_signed(-60, RAM(19)'LENGTH));
            ELSIF (number = 5) THEN
                RAM(8) <= STD_LOGIC_VECTOR(to_signed(20, RAM(19)'LENGTH));
                RAM(0) <= STD_LOGIC_VECTOR(to_signed(20, RAM(19)'LENGTH));
                RAM(18) <= STD_LOGIC_VECTOR(to_signed(20, RAM(19)'LENGTH));
                RAM(52) <= STD_LOGIC_VECTOR(to_signed(20, RAM(19)'LENGTH));
                RAM(64) <= STD_LOGIC_VECTOR(to_signed(-60, RAM(19)'LENGTH));
            ELSIF (number = 6) THEN
                RAM(8) <= STD_LOGIC_VECTOR(to_signed(20, RAM(19)'LENGTH));
                RAM(18) <= STD_LOGIC_VECTOR(to_signed(20, RAM(19)'LENGTH));
                RAM(57) <= STD_LOGIC_VECTOR(to_signed(20, RAM(19)'LENGTH));
                RAM(58) <= STD_LOGIC_VECTOR(to_signed(20, RAM(19)'LENGTH));
                RAM(67) <= STD_LOGIC_VECTOR(to_signed(-60, RAM(19)'LENGTH));
            ELSIF (number = 7) THEN
                RAM(9) <= STD_LOGIC_VECTOR(to_signed(20, RAM(19)'LENGTH));
                RAM(25) <= STD_LOGIC_VECTOR(to_signed(20, RAM(19)'LENGTH));
                RAM(27) <= STD_LOGIC_VECTOR(to_signed(20, RAM(19)'LENGTH));
                RAM(38) <= STD_LOGIC_VECTOR(to_signed(20, RAM(19)'LENGTH));
                RAM(65) <= STD_LOGIC_VECTOR(to_signed(-60, RAM(19)'LENGTH));
            ELSIF (number = 8) THEN
                RAM(12) <= STD_LOGIC_VECTOR(to_signed(20, RAM(19)'LENGTH));
                RAM(0) <= STD_LOGIC_VECTOR(to_signed(20, RAM(19)'LENGTH));
                RAM(20) <= STD_LOGIC_VECTOR(to_signed(20, RAM(19)'LENGTH));
                RAM(26) <= STD_LOGIC_VECTOR(to_signed(20, RAM(19)'LENGTH));
                RAM(63) <= STD_LOGIC_VECTOR(to_signed(-60, RAM(19)'LENGTH));
            ELSIF (number = 9) THEN
                RAM(15) <= STD_LOGIC_VECTOR(to_signed(20, RAM(19)'LENGTH));
                RAM(19) <= STD_LOGIC_VECTOR(to_signed(20, RAM(19)'LENGTH));
                RAM(47) <= STD_LOGIC_VECTOR(to_signed(20, RAM(19)'LENGTH));
                RAM(48) <= STD_LOGIC_VECTOR(to_signed(20, RAM(19)'LENGTH));
                RAM(65) <= STD_LOGIC_VECTOR(to_signed(-60, RAM(19)'LENGTH));
            ELSIF (number = 10) THEN
                RAM(8) <= STD_LOGIC_VECTOR(to_signed(20, RAM(19)'LENGTH));
                RAM(9) <= STD_LOGIC_VECTOR(to_signed(20, RAM(19)'LENGTH));
                RAM(18) <= STD_LOGIC_VECTOR(to_signed(20, RAM(19)'LENGTH));
                RAM(24) <= STD_LOGIC_VECTOR(to_signed(20, RAM(19)'LENGTH));
                RAM(65) <= STD_LOGIC_VECTOR(to_signed(-60, RAM(19)'LENGTH));
            ELSIF (number = 11) THEN
                RAM(15) <= STD_LOGIC_VECTOR(to_signed(20, RAM(19)'LENGTH));
                RAM(32) <= STD_LOGIC_VECTOR(to_signed(20, RAM(19)'LENGTH));
                RAM(35) <= STD_LOGIC_VECTOR(to_signed(20, RAM(19)'LENGTH));
                RAM(40) <= STD_LOGIC_VECTOR(to_signed(20, RAM(19)'LENGTH));
                RAM(62) <= STD_LOGIC_VECTOR(to_signed(-60, RAM(19)'LENGTH));
            ELSIF (number = 12) THEN
                RAM(2) <= STD_LOGIC_VECTOR(to_signed(20, RAM(19)'LENGTH));
                RAM(38) <= STD_LOGIC_VECTOR(to_signed(20, RAM(19)'LENGTH));
                RAM(41) <= STD_LOGIC_VECTOR(to_signed(20, RAM(19)'LENGTH));
                RAM(46) <= STD_LOGIC_VECTOR(to_signed(20, RAM(19)'LENGTH));
                RAM(63) <= STD_LOGIC_VECTOR(to_signed(-60, RAM(19)'LENGTH));
            ELSIF (number = 13) THEN
                RAM(7) <= STD_LOGIC_VECTOR(to_signed(20, RAM(19)'LENGTH));
                RAM(14) <= STD_LOGIC_VECTOR(to_signed(20, RAM(19)'LENGTH));
                RAM(0) <= STD_LOGIC_VECTOR(to_signed(20, RAM(19)'LENGTH));
                RAM(18) <= STD_LOGIC_VECTOR(to_signed(20, RAM(19)'LENGTH));
                RAM(70) <= STD_LOGIC_VECTOR(to_signed(-60, RAM(19)'LENGTH));
                RAM(0) <= STD_LOGIC_VECTOR(to_signed(4, RAM(19)'LENGTH));
            ELSIF (number = 14) THEN
                RAM(27) <= STD_LOGIC_VECTOR(to_signed(20, RAM(19)'LENGTH));
                RAM(37) <= STD_LOGIC_VECTOR(to_signed(20, RAM(19)'LENGTH));
                RAM(38) <= STD_LOGIC_VECTOR(to_signed(20, RAM(19)'LENGTH));
                RAM(49) <= STD_LOGIC_VECTOR(to_signed(20, RAM(19)'LENGTH));
                RAM(67) <= STD_LOGIC_VECTOR(to_signed(-60, RAM(19)'LENGTH));
            ELSIF (number = 15) THEN
                RAM(4) <= STD_LOGIC_VECTOR(to_signed(20, RAM(19)'LENGTH));
                RAM(34) <= STD_LOGIC_VECTOR(to_signed(20, RAM(19)'LENGTH));
                RAM(34) <= STD_LOGIC_VECTOR(to_signed(20, RAM(19)'LENGTH));
                RAM(35) <= STD_LOGIC_VECTOR(to_signed(20, RAM(19)'LENGTH));
                RAM(76) <= STD_LOGIC_VECTOR(to_signed(-60, RAM(19)'LENGTH));
            ELSIF (number = 16) THEN
                RAM(20) <= STD_LOGIC_VECTOR(to_signed(20, RAM(19)'LENGTH));
                RAM(20) <= STD_LOGIC_VECTOR(to_signed(20, RAM(19)'LENGTH));
                RAM(28) <= STD_LOGIC_VECTOR(to_signed(20, RAM(19)'LENGTH));
                RAM(61) <= STD_LOGIC_VECTOR(to_signed(20, RAM(19)'LENGTH));
                RAM(73) <= STD_LOGIC_VECTOR(to_signed(-60, RAM(19)'LENGTH));
            ELSIF (number = 17) THEN
                RAM(6) <= STD_LOGIC_VECTOR(to_signed(20, RAM(19)'LENGTH));
                RAM(35) <= STD_LOGIC_VECTOR(to_signed(20, RAM(19)'LENGTH));
                RAM(38) <= STD_LOGIC_VECTOR(to_signed(20, RAM(19)'LENGTH));
                RAM(40) <= STD_LOGIC_VECTOR(to_signed(20, RAM(19)'LENGTH));
                RAM(67) <= STD_LOGIC_VECTOR(to_signed(-60, RAM(19)'LENGTH));
            ELSIF (number = 18) THEN
                RAM(14) <= STD_LOGIC_VECTOR(to_signed(20, RAM(19)'LENGTH));
                RAM(23) <= STD_LOGIC_VECTOR(to_signed(20, RAM(19)'LENGTH));
                RAM(44) <= STD_LOGIC_VECTOR(to_signed(20, RAM(19)'LENGTH));
                RAM(49) <= STD_LOGIC_VECTOR(to_signed(20, RAM(19)'LENGTH));
                RAM(62) <= STD_LOGIC_VECTOR(to_signed(-60, RAM(19)'LENGTH));
            ELSIF (number = 19) THEN
                RAM(0) <= STD_LOGIC_VECTOR(to_signed(20, RAM(19)'LENGTH));
                RAM(18) <= STD_LOGIC_VECTOR(to_signed(20, RAM(19)'LENGTH));
                RAM(50) <= STD_LOGIC_VECTOR(to_signed(20, RAM(19)'LENGTH));
                RAM(53) <= STD_LOGIC_VECTOR(to_signed(20, RAM(19)'LENGTH));
                RAM(63) <= STD_LOGIC_VECTOR(to_signed(-60, RAM(19)'LENGTH));
            ELSIF (number = 20) THEN
                RAM(7) <= STD_LOGIC_VECTOR(to_signed(20, RAM(19)'LENGTH));
                RAM(22) <= STD_LOGIC_VECTOR(to_signed(20, RAM(19)'LENGTH));
                RAM(31) <= STD_LOGIC_VECTOR(to_signed(20, RAM(19)'LENGTH));
                RAM(59) <= STD_LOGIC_VECTOR(to_signed(20, RAM(19)'LENGTH));
                RAM(62) <= STD_LOGIC_VECTOR(to_signed(-60, RAM(19)'LENGTH));
            ELSIF (number = 21) THEN
                RAM(0) <= STD_LOGIC_VECTOR(to_signed(20, RAM(19)'LENGTH));
                RAM(23) <= STD_LOGIC_VECTOR(to_signed(20, RAM(19)'LENGTH));
                RAM(48) <= STD_LOGIC_VECTOR(to_signed(20, RAM(19)'LENGTH));
                RAM(52) <= STD_LOGIC_VECTOR(to_signed(20, RAM(19)'LENGTH));
                RAM(68) <= STD_LOGIC_VECTOR(to_signed(-60, RAM(19)'LENGTH));
            ELSIF (number = 22) THEN
                RAM(7) <= STD_LOGIC_VECTOR(to_signed(20, RAM(19)'LENGTH));
                RAM(19) <= STD_LOGIC_VECTOR(to_signed(20, RAM(19)'LENGTH));
                RAM(21) <= STD_LOGIC_VECTOR(to_signed(20, RAM(19)'LENGTH));
                RAM(22) <= STD_LOGIC_VECTOR(to_signed(20, RAM(19)'LENGTH));
                RAM(69) <= STD_LOGIC_VECTOR(to_signed(-60, RAM(19)'LENGTH));
            ELSIF (number = 23) THEN
                RAM(9) <= STD_LOGIC_VECTOR(to_signed(20, RAM(19)'LENGTH));
                RAM(20) <= STD_LOGIC_VECTOR(to_signed(20, RAM(19)'LENGTH));
                RAM(11) <= STD_LOGIC_VECTOR(to_signed(20, RAM(19)'LENGTH));
                RAM(30) <= STD_LOGIC_VECTOR(to_signed(20, RAM(19)'LENGTH));
                RAM(67) <= STD_LOGIC_VECTOR(to_signed(-60, RAM(19)'LENGTH));
            ELSIF (number = 24) THEN
                RAM(14) <= STD_LOGIC_VECTOR(to_signed(20, RAM(19)'LENGTH));
                RAM(19) <= STD_LOGIC_VECTOR(to_signed(20, RAM(19)'LENGTH));
                RAM(43) <= STD_LOGIC_VECTOR(to_signed(20, RAM(19)'LENGTH));
                RAM(59) <= STD_LOGIC_VECTOR(to_signed(20, RAM(19)'LENGTH));
                RAM(76) <= STD_LOGIC_VECTOR(to_signed(-60, RAM(19)'LENGTH));
            ELSIF (number = 25) THEN
                RAM(25) <= STD_LOGIC_VECTOR(to_signed(20, RAM(19)'LENGTH));
                RAM(30) <= STD_LOGIC_VECTOR(to_signed(20, RAM(19)'LENGTH));
                RAM(33) <= STD_LOGIC_VECTOR(to_signed(20, RAM(19)'LENGTH));
                RAM(48) <= STD_LOGIC_VECTOR(to_signed(20, RAM(19)'LENGTH));
                RAM(74) <= STD_LOGIC_VECTOR(to_signed(-60, RAM(19)'LENGTH));
            ELSIF (number = 26) THEN
                RAM(18) <= STD_LOGIC_VECTOR(to_signed(20, RAM(19)'LENGTH));
                RAM(31) <= STD_LOGIC_VECTOR(to_signed(20, RAM(19)'LENGTH));
                RAM(32) <= STD_LOGIC_VECTOR(to_signed(20, RAM(19)'LENGTH));
                RAM(42) <= STD_LOGIC_VECTOR(to_signed(20, RAM(19)'LENGTH));
                RAM(65) <= STD_LOGIC_VECTOR(to_signed(-60, RAM(19)'LENGTH));
            ELSIF (number = 27) THEN
                RAM(20) <= STD_LOGIC_VECTOR(to_signed(20, RAM(19)'LENGTH));
                RAM(15) <= STD_LOGIC_VECTOR(to_signed(20, RAM(19)'LENGTH));
                RAM(49) <= STD_LOGIC_VECTOR(to_signed(20, RAM(19)'LENGTH));
                RAM(51) <= STD_LOGIC_VECTOR(to_signed(20, RAM(19)'LENGTH));
                RAM(75) <= STD_LOGIC_VECTOR(to_signed(-60, RAM(19)'LENGTH));
            ELSIF (number = 28) THEN
                RAM(3) <= STD_LOGIC_VECTOR(to_signed(20, RAM(19)'LENGTH));
                RAM(40) <= STD_LOGIC_VECTOR(to_signed(20, RAM(19)'LENGTH));
                RAM(51) <= STD_LOGIC_VECTOR(to_signed(20, RAM(19)'LENGTH));
                RAM(52) <= STD_LOGIC_VECTOR(to_signed(20, RAM(19)'LENGTH));
                RAM(65) <= STD_LOGIC_VECTOR(to_signed(-60, RAM(19)'LENGTH));
            ELSIF (number = 29) THEN
                RAM(7) <= STD_LOGIC_VECTOR(to_signed(20, RAM(19)'LENGTH));
                RAM(8) <= STD_LOGIC_VECTOR(to_signed(20, RAM(19)'LENGTH));
                RAM(20) <= STD_LOGIC_VECTOR(to_signed(20, RAM(19)'LENGTH));
                RAM(30) <= STD_LOGIC_VECTOR(to_signed(20, RAM(19)'LENGTH));
                RAM(64) <= STD_LOGIC_VECTOR(to_signed(-60, RAM(19)'LENGTH));
            ELSIF (number = 30) THEN
                RAM(11) <= STD_LOGIC_VECTOR(to_signed(20, RAM(19)'LENGTH));
                RAM(12) <= STD_LOGIC_VECTOR(to_signed(20, RAM(19)'LENGTH));
                RAM(18) <= STD_LOGIC_VECTOR(to_signed(20, RAM(19)'LENGTH));
                RAM(39) <= STD_LOGIC_VECTOR(to_signed(20, RAM(19)'LENGTH));
                RAM(65) <= STD_LOGIC_VECTOR(to_signed(-60, RAM(19)'LENGTH));
            ELSIF (number = 31) THEN
                RAM(8) <= STD_LOGIC_VECTOR(to_signed(20, RAM(19)'LENGTH));
                RAM(18) <= STD_LOGIC_VECTOR(to_signed(20, RAM(19)'LENGTH));
                RAM(55) <= STD_LOGIC_VECTOR(to_signed(20, RAM(19)'LENGTH));
                RAM(59) <= STD_LOGIC_VECTOR(to_signed(20, RAM(19)'LENGTH));
                RAM(72) <= STD_LOGIC_VECTOR(to_signed(-60, RAM(19)'LENGTH));
            ELSIF (number = 32) THEN
                RAM(9) <= STD_LOGIC_VECTOR(to_signed(20, RAM(19)'LENGTH));
                RAM(14) <= STD_LOGIC_VECTOR(to_signed(20, RAM(19)'LENGTH));
                RAM(23) <= STD_LOGIC_VECTOR(to_signed(20, RAM(19)'LENGTH));
                RAM(50) <= STD_LOGIC_VECTOR(to_signed(20, RAM(19)'LENGTH));
                RAM(65) <= STD_LOGIC_VECTOR(to_signed(-60, RAM(19)'LENGTH));
            ELSIF (number = 33) THEN
                RAM(2) <= STD_LOGIC_VECTOR(to_signed(20, RAM(19)'LENGTH));
                RAM(18) <= STD_LOGIC_VECTOR(to_signed(20, RAM(19)'LENGTH));
                RAM(19) <= STD_LOGIC_VECTOR(to_signed(20, RAM(19)'LENGTH));
                RAM(47) <= STD_LOGIC_VECTOR(to_signed(20, RAM(19)'LENGTH));
                RAM(68) <= STD_LOGIC_VECTOR(to_signed(-60, RAM(19)'LENGTH));
            ELSIF (number = 34) THEN
                RAM(8) <= STD_LOGIC_VECTOR(to_signed(20, RAM(19)'LENGTH));
                RAM(14) <= STD_LOGIC_VECTOR(to_signed(20, RAM(19)'LENGTH));
                RAM(31) <= STD_LOGIC_VECTOR(to_signed(20, RAM(19)'LENGTH));
                RAM(33) <= STD_LOGIC_VECTOR(to_signed(20, RAM(19)'LENGTH));
                RAM(65) <= STD_LOGIC_VECTOR(to_signed(-60, RAM(19)'LENGTH));
            ELSIF (number = 35) THEN
                RAM(0) <= STD_LOGIC_VECTOR(to_signed(20, RAM(19)'LENGTH));
                RAM(26) <= STD_LOGIC_VECTOR(to_signed(20, RAM(19)'LENGTH));
                RAM(55) <= STD_LOGIC_VECTOR(to_signed(20, RAM(19)'LENGTH));
                RAM(60) <= STD_LOGIC_VECTOR(to_signed(20, RAM(19)'LENGTH));
                RAM(72) <= STD_LOGIC_VECTOR(to_signed(-60, RAM(19)'LENGTH));
            ELSIF (number = 36) THEN
                RAM(13) <= STD_LOGIC_VECTOR(to_signed(20, RAM(19)'LENGTH));
                RAM(30) <= STD_LOGIC_VECTOR(to_signed(20, RAM(19)'LENGTH));
                RAM(42) <= STD_LOGIC_VECTOR(to_signed(20, RAM(19)'LENGTH));
                RAM(51) <= STD_LOGIC_VECTOR(to_signed(20, RAM(19)'LENGTH));
                RAM(70) <= STD_LOGIC_VECTOR(to_signed(-60, RAM(19)'LENGTH));
            ELSIF (number = 37) THEN
                RAM(4) <= STD_LOGIC_VECTOR(to_signed(20, RAM(19)'LENGTH));
                RAM(15) <= STD_LOGIC_VECTOR(to_signed(20, RAM(19)'LENGTH));
                RAM(39) <= STD_LOGIC_VECTOR(to_signed(20, RAM(19)'LENGTH));
                RAM(58) <= STD_LOGIC_VECTOR(to_signed(20, RAM(19)'LENGTH));
                RAM(64) <= STD_LOGIC_VECTOR(to_signed(-60, RAM(19)'LENGTH));
            ELSIF (number = 38) THEN
                RAM(13) <= STD_LOGIC_VECTOR(to_signed(20, RAM(19)'LENGTH));
                RAM(18) <= STD_LOGIC_VECTOR(to_signed(20, RAM(19)'LENGTH));
                RAM(34) <= STD_LOGIC_VECTOR(to_signed(20, RAM(19)'LENGTH));
                RAM(55) <= STD_LOGIC_VECTOR(to_signed(20, RAM(19)'LENGTH));
                RAM(63) <= STD_LOGIC_VECTOR(to_signed(-60, RAM(19)'LENGTH));
            ELSIF (number = 39) THEN
                RAM(7) <= STD_LOGIC_VECTOR(to_signed(20, RAM(19)'LENGTH));
                RAM(19) <= STD_LOGIC_VECTOR(to_signed(20, RAM(19)'LENGTH));
                RAM(27) <= STD_LOGIC_VECTOR(to_signed(20, RAM(19)'LENGTH));
                RAM(30) <= STD_LOGIC_VECTOR(to_signed(20, RAM(19)'LENGTH));
                RAM(73) <= STD_LOGIC_VECTOR(to_signed(-60, RAM(19)'LENGTH));
            ELSIF (number = 40) THEN
                RAM(14) <= STD_LOGIC_VECTOR(to_signed(20, RAM(19)'LENGTH));
                RAM(27) <= STD_LOGIC_VECTOR(to_signed(20, RAM(19)'LENGTH));
                RAM(30) <= STD_LOGIC_VECTOR(to_signed(20, RAM(19)'LENGTH));
                RAM(34) <= STD_LOGIC_VECTOR(to_signed(20, RAM(19)'LENGTH));
                RAM(65) <= STD_LOGIC_VECTOR(to_signed(-60, RAM(19)'LENGTH));
            ELSIF (number = 41) THEN
                RAM(5) <= STD_LOGIC_VECTOR(to_signed(20, RAM(19)'LENGTH));
                RAM(14) <= STD_LOGIC_VECTOR(to_signed(20, RAM(19)'LENGTH));
                RAM(43) <= STD_LOGIC_VECTOR(to_signed(20, RAM(19)'LENGTH));
                RAM(57) <= STD_LOGIC_VECTOR(to_signed(20, RAM(19)'LENGTH));
                RAM(67) <= STD_LOGIC_VECTOR(to_signed(-60, RAM(19)'LENGTH));
            ELSIF (number = 42) THEN
                RAM(0) <= STD_LOGIC_VECTOR(to_signed(20, RAM(19)'LENGTH));
                RAM(34) <= STD_LOGIC_VECTOR(to_signed(20, RAM(19)'LENGTH));
                RAM(43) <= STD_LOGIC_VECTOR(to_signed(20, RAM(19)'LENGTH));
                RAM(45) <= STD_LOGIC_VECTOR(to_signed(20, RAM(19)'LENGTH));
                RAM(67) <= STD_LOGIC_VECTOR(to_signed(-60, RAM(19)'LENGTH));
            ELSIF (number = 43) THEN
                RAM(18) <= STD_LOGIC_VECTOR(to_signed(20, RAM(19)'LENGTH));
                RAM(29) <= STD_LOGIC_VECTOR(to_signed(20, RAM(19)'LENGTH));
                RAM(38) <= STD_LOGIC_VECTOR(to_signed(20, RAM(19)'LENGTH));
                RAM(53) <= STD_LOGIC_VECTOR(to_signed(20, RAM(19)'LENGTH));
                RAM(69) <= STD_LOGIC_VECTOR(to_signed(-60, RAM(19)'LENGTH));
            ELSIF (number = 44) THEN
                RAM(23) <= STD_LOGIC_VECTOR(to_signed(20, RAM(19)'LENGTH));
                RAM(25) <= STD_LOGIC_VECTOR(to_signed(20, RAM(19)'LENGTH));
                RAM(47) <= STD_LOGIC_VECTOR(to_signed(20, RAM(19)'LENGTH));
                RAM(50) <= STD_LOGIC_VECTOR(to_signed(20, RAM(19)'LENGTH));
                RAM(68) <= STD_LOGIC_VECTOR(to_signed(-60, RAM(19)'LENGTH));
            ELSIF (number = 45) THEN
                RAM(9) <= STD_LOGIC_VECTOR(to_signed(20, RAM(19)'LENGTH));
                RAM(12) <= STD_LOGIC_VECTOR(to_signed(20, RAM(19)'LENGTH));
                RAM(20) <= STD_LOGIC_VECTOR(to_signed(20, RAM(19)'LENGTH));
                RAM(36) <= STD_LOGIC_VECTOR(to_signed(20, RAM(19)'LENGTH));
                RAM(65) <= STD_LOGIC_VECTOR(to_signed(-60, RAM(19)'LENGTH));
            ELSIF (number = 46) THEN
                RAM(27) <= STD_LOGIC_VECTOR(to_signed(20, RAM(19)'LENGTH));
                RAM(33) <= STD_LOGIC_VECTOR(to_signed(20, RAM(19)'LENGTH));
                RAM(51) <= STD_LOGIC_VECTOR(to_signed(20, RAM(19)'LENGTH));
                RAM(52) <= STD_LOGIC_VECTOR(to_signed(20, RAM(19)'LENGTH));
                RAM(74) <= STD_LOGIC_VECTOR(to_signed(-60, RAM(19)'LENGTH));
            ELSIF (number = 47) THEN
                RAM(19) <= STD_LOGIC_VECTOR(to_signed(20, RAM(19)'LENGTH));
                RAM(27) <= STD_LOGIC_VECTOR(to_signed(20, RAM(19)'LENGTH));
                RAM(33) <= STD_LOGIC_VECTOR(to_signed(20, RAM(19)'LENGTH));
                RAM(56) <= STD_LOGIC_VECTOR(to_signed(20, RAM(19)'LENGTH));
                RAM(68) <= STD_LOGIC_VECTOR(to_signed(-60, RAM(19)'LENGTH));
            ELSIF (number = 48) THEN
                RAM(20) <= STD_LOGIC_VECTOR(to_signed(20, RAM(19)'LENGTH));
                RAM(18) <= STD_LOGIC_VECTOR(to_signed(20, RAM(19)'LENGTH));
                RAM(19) <= STD_LOGIC_VECTOR(to_signed(20, RAM(19)'LENGTH));
                RAM(49) <= STD_LOGIC_VECTOR(to_signed(20, RAM(19)'LENGTH));
                RAM(72) <= STD_LOGIC_VECTOR(to_signed(-60, RAM(19)'LENGTH));
            ELSIF (number = 49) THEN
                RAM(8) <= STD_LOGIC_VECTOR(to_signed(20, RAM(19)'LENGTH));
                RAM(12) <= STD_LOGIC_VECTOR(to_signed(20, RAM(19)'LENGTH));
                RAM(14) <= STD_LOGIC_VECTOR(to_signed(20, RAM(19)'LENGTH));
                RAM(57) <= STD_LOGIC_VECTOR(to_signed(20, RAM(19)'LENGTH));
                RAM(74) <= STD_LOGIC_VECTOR(to_signed(-60, RAM(19)'LENGTH));
            ELSIF (number = 50) THEN
                RAM(31) <= STD_LOGIC_VECTOR(to_signed(20, RAM(19)'LENGTH));
                RAM(52) <= STD_LOGIC_VECTOR(to_signed(20, RAM(19)'LENGTH));
                RAM(55) <= STD_LOGIC_VECTOR(to_signed(20, RAM(19)'LENGTH));
                RAM(59) <= STD_LOGIC_VECTOR(to_signed(20, RAM(19)'LENGTH));
                RAM(73) <= STD_LOGIC_VECTOR(to_signed(-60, RAM(19)'LENGTH));
            ELSIF (number = 51) THEN
                RAM(7) <= STD_LOGIC_VECTOR(to_signed(20, RAM(19)'LENGTH));
                RAM(20) <= STD_LOGIC_VECTOR(to_signed(20, RAM(19)'LENGTH));
                RAM(16) <= STD_LOGIC_VECTOR(to_signed(20, RAM(19)'LENGTH));
                RAM(0) <= STD_LOGIC_VECTOR(to_signed(20, RAM(19)'LENGTH));
                RAM(68) <= STD_LOGIC_VECTOR(to_signed(-60, RAM(19)'LENGTH));
            ELSIF (number = 52) THEN
                RAM(2) <= STD_LOGIC_VECTOR(to_signed(20, RAM(19)'LENGTH));
                RAM(27) <= STD_LOGIC_VECTOR(to_signed(20, RAM(19)'LENGTH));
                RAM(53) <= STD_LOGIC_VECTOR(to_signed(20, RAM(19)'LENGTH));
                RAM(58) <= STD_LOGIC_VECTOR(to_signed(20, RAM(19)'LENGTH));
                RAM(69) <= STD_LOGIC_VECTOR(to_signed(-60, RAM(19)'LENGTH));
            ELSIF (number = 53) THEN
                RAM(2) <= STD_LOGIC_VECTOR(to_signed(20, RAM(19)'LENGTH));
                RAM(21) <= STD_LOGIC_VECTOR(to_signed(20, RAM(19)'LENGTH));
                RAM(36) <= STD_LOGIC_VECTOR(to_signed(20, RAM(19)'LENGTH));
                RAM(47) <= STD_LOGIC_VECTOR(to_signed(20, RAM(19)'LENGTH));
                RAM(71) <= STD_LOGIC_VECTOR(to_signed(-60, RAM(19)'LENGTH));
            ELSIF (number = 54) THEN
                RAM(32) <= STD_LOGIC_VECTOR(to_signed(20, RAM(19)'LENGTH));
                RAM(34) <= STD_LOGIC_VECTOR(to_signed(20, RAM(19)'LENGTH));
                RAM(48) <= STD_LOGIC_VECTOR(to_signed(20, RAM(19)'LENGTH));
                RAM(56) <= STD_LOGIC_VECTOR(to_signed(20, RAM(19)'LENGTH));
                RAM(70) <= STD_LOGIC_VECTOR(to_signed(-60, RAM(19)'LENGTH));
            ELSIF (number = 55) THEN
                RAM(7) <= STD_LOGIC_VECTOR(to_signed(20, RAM(19)'LENGTH));
                RAM(42) <= STD_LOGIC_VECTOR(to_signed(20, RAM(19)'LENGTH));
                RAM(50) <= STD_LOGIC_VECTOR(to_signed(20, RAM(19)'LENGTH));
                RAM(52) <= STD_LOGIC_VECTOR(to_signed(20, RAM(19)'LENGTH));
                RAM(70) <= STD_LOGIC_VECTOR(to_signed(-60, RAM(19)'LENGTH));
            ELSIF (number = 56) THEN
                RAM(12) <= STD_LOGIC_VECTOR(to_signed(20, RAM(19)'LENGTH));
                RAM(12) <= STD_LOGIC_VECTOR(to_signed(20, RAM(19)'LENGTH));
                RAM(27) <= STD_LOGIC_VECTOR(to_signed(20, RAM(19)'LENGTH));
                RAM(37) <= STD_LOGIC_VECTOR(to_signed(20, RAM(19)'LENGTH));
                RAM(68) <= STD_LOGIC_VECTOR(to_signed(-60, RAM(19)'LENGTH));
            ELSIF (number = 57) THEN
                RAM(40) <= STD_LOGIC_VECTOR(to_signed(20, RAM(19)'LENGTH));
                RAM(40) <= STD_LOGIC_VECTOR(to_signed(20, RAM(19)'LENGTH));
                RAM(41) <= STD_LOGIC_VECTOR(to_signed(20, RAM(19)'LENGTH));
                RAM(59) <= STD_LOGIC_VECTOR(to_signed(20, RAM(19)'LENGTH));
                RAM(67) <= STD_LOGIC_VECTOR(to_signed(-60, RAM(19)'LENGTH));
            ELSIF (number = 58) THEN
                RAM(20) <= STD_LOGIC_VECTOR(to_signed(20, RAM(19)'LENGTH));
                RAM(34) <= STD_LOGIC_VECTOR(to_signed(20, RAM(19)'LENGTH));
                RAM(44) <= STD_LOGIC_VECTOR(to_signed(20, RAM(19)'LENGTH));
                RAM(49) <= STD_LOGIC_VECTOR(to_signed(20, RAM(19)'LENGTH));
                RAM(72) <= STD_LOGIC_VECTOR(to_signed(-60, RAM(19)'LENGTH));
            ELSIF (number = 59) THEN
                RAM(25) <= STD_LOGIC_VECTOR(to_signed(20, RAM(19)'LENGTH));
                RAM(29) <= STD_LOGIC_VECTOR(to_signed(20, RAM(19)'LENGTH));
                RAM(41) <= STD_LOGIC_VECTOR(to_signed(20, RAM(19)'LENGTH));
                RAM(59) <= STD_LOGIC_VECTOR(to_signed(20, RAM(19)'LENGTH));
                RAM(62) <= STD_LOGIC_VECTOR(to_signed(-60, RAM(19)'LENGTH));
            ELSIF (number = 60) THEN
                RAM(25) <= STD_LOGIC_VECTOR(to_signed(20, RAM(19)'LENGTH));
                RAM(46) <= STD_LOGIC_VECTOR(to_signed(20, RAM(19)'LENGTH));
                RAM(47) <= STD_LOGIC_VECTOR(to_signed(20, RAM(19)'LENGTH));
                RAM(47) <= STD_LOGIC_VECTOR(to_signed(20, RAM(19)'LENGTH));
                RAM(64) <= STD_LOGIC_VECTOR(to_signed(-60, RAM(19)'LENGTH));
            ELSIF (number = 61) THEN
                RAM(2) <= STD_LOGIC_VECTOR(to_signed(20, RAM(19)'LENGTH));
                RAM(20) <= STD_LOGIC_VECTOR(to_signed(20, RAM(19)'LENGTH));
                RAM(15) <= STD_LOGIC_VECTOR(to_signed(20, RAM(19)'LENGTH));
                RAM(39) <= STD_LOGIC_VECTOR(to_signed(20, RAM(19)'LENGTH));
                RAM(68) <= STD_LOGIC_VECTOR(to_signed(-60, RAM(19)'LENGTH));
            ELSIF (number = 62) THEN
                RAM(9) <= STD_LOGIC_VECTOR(to_signed(85, RAM(19)'LENGTH));
                RAM(33) <= STD_LOGIC_VECTOR(to_signed(85, RAM(19)'LENGTH));
                RAM(38) <= STD_LOGIC_VECTOR(to_signed(85, RAM(19)'LENGTH));
                RAM(38) <= STD_LOGIC_VECTOR(to_signed(85, RAM(19)'LENGTH));
                RAM(63) <= STD_LOGIC_VECTOR(to_signed(-60, RAM(19)'LENGTH));
            ELSIF (number = 63) THEN
                RAM(19) <= STD_LOGIC_VECTOR(to_signed(85, RAM(19)'LENGTH));
                RAM(22) <= STD_LOGIC_VECTOR(to_signed(85, RAM(19)'LENGTH));
                RAM(36) <= STD_LOGIC_VECTOR(to_signed(85, RAM(19)'LENGTH));
                RAM(52) <= STD_LOGIC_VECTOR(to_signed(85, RAM(19)'LENGTH));
                RAM(68) <= STD_LOGIC_VECTOR(to_signed(-60, RAM(19)'LENGTH));
            ELSIF (number = 64) THEN
                RAM(18) <= STD_LOGIC_VECTOR(to_signed(85, RAM(19)'LENGTH));
                RAM(23) <= STD_LOGIC_VECTOR(to_signed(85, RAM(19)'LENGTH));
                RAM(23) <= STD_LOGIC_VECTOR(to_signed(85, RAM(19)'LENGTH));
                RAM(24) <= STD_LOGIC_VECTOR(to_signed(85, RAM(19)'LENGTH));
                RAM(64) <= STD_LOGIC_VECTOR(to_signed(-60, RAM(19)'LENGTH));
            ELSIF (number = 65) THEN
                RAM(4) <= STD_LOGIC_VECTOR(to_signed(85, RAM(19)'LENGTH));
                RAM(32) <= STD_LOGIC_VECTOR(to_signed(85, RAM(19)'LENGTH));
                RAM(38) <= STD_LOGIC_VECTOR(to_signed(85, RAM(19)'LENGTH));
                RAM(40) <= STD_LOGIC_VECTOR(to_signed(85, RAM(19)'LENGTH));
                RAM(62) <= STD_LOGIC_VECTOR(to_signed(-60, RAM(19)'LENGTH));
            ELSIF (number = 66) THEN
                RAM(2) <= STD_LOGIC_VECTOR(to_signed(85, RAM(19)'LENGTH));
                RAM(20) <= STD_LOGIC_VECTOR(to_signed(85, RAM(19)'LENGTH));
                RAM(26) <= STD_LOGIC_VECTOR(to_signed(85, RAM(19)'LENGTH));
                RAM(59) <= STD_LOGIC_VECTOR(to_signed(85, RAM(19)'LENGTH));
                RAM(71) <= STD_LOGIC_VECTOR(to_signed(-60, RAM(19)'LENGTH));
            ELSIF (number = 67) THEN
                RAM(20) <= STD_LOGIC_VECTOR(to_signed(85, RAM(19)'LENGTH));
                RAM(40) <= STD_LOGIC_VECTOR(to_signed(85, RAM(19)'LENGTH));
                RAM(44) <= STD_LOGIC_VECTOR(to_signed(85, RAM(19)'LENGTH));
                RAM(48) <= STD_LOGIC_VECTOR(to_signed(85, RAM(19)'LENGTH));
                RAM(63) <= STD_LOGIC_VECTOR(to_signed(-60, RAM(19)'LENGTH));
            ELSIF (number = 68) THEN
                RAM(20) <= STD_LOGIC_VECTOR(to_signed(85, RAM(19)'LENGTH));
                RAM(15) <= STD_LOGIC_VECTOR(to_signed(85, RAM(19)'LENGTH));
                RAM(42) <= STD_LOGIC_VECTOR(to_signed(85, RAM(19)'LENGTH));
                RAM(50) <= STD_LOGIC_VECTOR(to_signed(85, RAM(19)'LENGTH));
                RAM(69) <= STD_LOGIC_VECTOR(to_signed(-60, RAM(19)'LENGTH));
            ELSIF (number = 69) THEN
                RAM(25) <= STD_LOGIC_VECTOR(to_signed(85, RAM(19)'LENGTH));
                RAM(25) <= STD_LOGIC_VECTOR(to_signed(85, RAM(19)'LENGTH));
                RAM(34) <= STD_LOGIC_VECTOR(to_signed(85, RAM(19)'LENGTH));
                RAM(46) <= STD_LOGIC_VECTOR(to_signed(85, RAM(19)'LENGTH));
                RAM(69) <= STD_LOGIC_VECTOR(to_signed(-60, RAM(19)'LENGTH));
            ELSIF (number = 70) THEN
                RAM(13) <= STD_LOGIC_VECTOR(to_signed(85, RAM(19)'LENGTH));
                RAM(24) <= STD_LOGIC_VECTOR(to_signed(85, RAM(19)'LENGTH));
                RAM(32) <= STD_LOGIC_VECTOR(to_signed(85, RAM(19)'LENGTH));
                RAM(50) <= STD_LOGIC_VECTOR(to_signed(85, RAM(19)'LENGTH));
                RAM(63) <= STD_LOGIC_VECTOR(to_signed(-60, RAM(19)'LENGTH));
            ELSIF (number = 71) THEN
                RAM(5) <= STD_LOGIC_VECTOR(to_signed(85, RAM(19)'LENGTH));
                RAM(32) <= STD_LOGIC_VECTOR(to_signed(85, RAM(19)'LENGTH));
                RAM(60) <= STD_LOGIC_VECTOR(to_signed(85, RAM(19)'LENGTH));
                RAM(61) <= STD_LOGIC_VECTOR(to_signed(85, RAM(19)'LENGTH));
                RAM(65) <= STD_LOGIC_VECTOR(to_signed(-60, RAM(19)'LENGTH));
                RAM(1) <= STD_LOGIC_VECTOR(to_signed(4, RAM(19)'LENGTH));
            ELSIF (number = 72) THEN
                RAM(15) <= STD_LOGIC_VECTOR(to_signed(85, RAM(19)'LENGTH));
                RAM(27) <= STD_LOGIC_VECTOR(to_signed(85, RAM(19)'LENGTH));
                RAM(33) <= STD_LOGIC_VECTOR(to_signed(85, RAM(19)'LENGTH));
                RAM(48) <= STD_LOGIC_VECTOR(to_signed(85, RAM(19)'LENGTH));
                RAM(67) <= STD_LOGIC_VECTOR(to_signed(-60, RAM(19)'LENGTH));
            ELSIF (number = 73) THEN
                RAM(3) <= STD_LOGIC_VECTOR(to_signed(85, RAM(19)'LENGTH));
                RAM(28) <= STD_LOGIC_VECTOR(to_signed(85, RAM(19)'LENGTH));
                RAM(48) <= STD_LOGIC_VECTOR(to_signed(85, RAM(19)'LENGTH));
                RAM(50) <= STD_LOGIC_VECTOR(to_signed(85, RAM(19)'LENGTH));
                RAM(72) <= STD_LOGIC_VECTOR(to_signed(-60, RAM(19)'LENGTH));
            ELSIF (number = 74) THEN
                RAM(12) <= STD_LOGIC_VECTOR(to_signed(85, RAM(19)'LENGTH));
                RAM(45) <= STD_LOGIC_VECTOR(to_signed(85, RAM(19)'LENGTH));
                RAM(47) <= STD_LOGIC_VECTOR(to_signed(85, RAM(19)'LENGTH));
                RAM(53) <= STD_LOGIC_VECTOR(to_signed(85, RAM(19)'LENGTH));
                RAM(70) <= STD_LOGIC_VECTOR(to_signed(-60, RAM(19)'LENGTH));
            ELSIF (number = 75) THEN
                RAM(2) <= STD_LOGIC_VECTOR(to_signed(85, RAM(19)'LENGTH));
                RAM(13) <= STD_LOGIC_VECTOR(to_signed(85, RAM(19)'LENGTH));
                RAM(47) <= STD_LOGIC_VECTOR(to_signed(85, RAM(19)'LENGTH));
                RAM(54) <= STD_LOGIC_VECTOR(to_signed(85, RAM(19)'LENGTH));
                RAM(71) <= STD_LOGIC_VECTOR(to_signed(-60, RAM(19)'LENGTH));
            ELSIF (number = 76) THEN
                RAM(12) <= STD_LOGIC_VECTOR(to_signed(85, RAM(19)'LENGTH));
                RAM(25) <= STD_LOGIC_VECTOR(to_signed(85, RAM(19)'LENGTH));
                RAM(44) <= STD_LOGIC_VECTOR(to_signed(85, RAM(19)'LENGTH));
                RAM(61) <= STD_LOGIC_VECTOR(to_signed(85, RAM(19)'LENGTH));
                RAM(62) <= STD_LOGIC_VECTOR(to_signed(-60, RAM(19)'LENGTH));

            END IF;
        END IF;
        IF dpra = x"ff" THEN
            dpo <= STD_LOGIC_VECTOR(to_signed(20, RAM(19)'LENGTH));
        ELSE
            dpo <= RAM(conv_integer(dpra));
        END IF;
    END PROCESS;
END syn;